`timescale 1ns/1ns
`include "head.v"
module ALU (
	input [2:0] ALUCtrl,
    input [31:0] A,
    input [31:0] B,
    output [31:0] C
    );


wire [31:0] out = (A[31] == 1) ? 0:
                  (A[30] == 1) ? 1:
                  (A[29] == 1) ? 2:
                  (A[28] == 1) ? 3:
                  (A[27] == 1) ? 4:
                  (A[26] == 1) ? 5:
                  (A[25] == 1) ? 6:
                  (A[24] == 1) ? 7:
                  (A[23] == 1) ? 8:
                  (A[22] == 1) ? 9:
                  (A[21] == 1) ? 10:
                  (A[20] == 1) ? 11:
                  (A[19] == 1) ? 12:
                  (A[18] == 1) ? 13:
                  (A[17] == 1) ? 14:
                  (A[16] == 1) ? 15:
                  (A[15] == 1) ? 16:
                  (A[14] == 1) ? 17:
                  (A[13] == 1) ? 18:
                  (A[12] == 1) ? 19:
                  (A[11] == 1) ? 20:
                  (A[10] == 1) ? 21:
                   (A[9] == 1) ? 22:
                   (A[8] == 1) ? 23:
                   (A[7] == 1) ? 24:
                   (A[6] == 1) ? 25:
                   (A[5] == 1) ? 26:
                   (A[4] == 1) ? 27:
                   (A[3] == 1) ? 28:
                   (A[2] == 1) ? 29:
                   (A[1] == 1) ? 30:
                   (A[0] == 1) ? 31:
                                 32;

	assign C = (ALUCtrl == `ALU_SUBU) ? A - B:
				 (ALUCtrl == `ALU_OR) ? A | B:
				 (ALUCtrl == `ALU_CLZ) ? out:
									   A + B;


    
endmodule